
package test_pkg;
  import uvm_pkg::*;
 `include "monitor.svh"

endpackage


