`timescale 1ns / 1ns


interface dut_if;

    reg  clk;
    reg[7:0] in;
    reg rst;
    wire  out; 
    reg [7:0] in_last;

endinterface



    
    




